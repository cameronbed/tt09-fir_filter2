//------> /eda/mentor/Siemens_EDA/Catapult_Synthesis_2023.1_2/Mgc_home/pkgs/siflibs/ccs_out_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

module ccs_out_v1 (dat, idat);

  // parameter integer rscid = 1;
  parameter integer width = 8;

  output   [width-1:0] dat;
  input    [width-1:0] idat;

  wire     [width-1:0] dat;

  assign dat = idat;

endmodule




//------> /eda/mentor/Siemens_EDA/Catapult_Synthesis_2023.1_2/Mgc_home/pkgs/siflibs/ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_in_v1 (idat, dat);

  // 
  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> /eda/mentor/Siemens_EDA/Catapult_Synthesis_2023.1_2/Mgc_home/pkgs/siflibs/mgc_io_sync_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module mgc_io_sync_v2 (ld, lz);
    parameter valid = 0;

    input  ld;
    output lz;

    wire   lz;

    assign lz = ld;

endmodule


//------> ./rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2023.1_2/1049935 Production Release
//  HLS Date:       Sat Jun 10 10:53:51 PDT 2023
// 
//  Generated by:   hx2227@hansolo.poly.edu
//  Generated date: Wed Dec 11 13:34:35 2024
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    fir_core_core_fsm
//  FSM Module
// ------------------------------------------------------------------


module fir_core_core_fsm (
  clk, rst, fsm_output, Shift_Accum_Loop_C_5_tr0
);
  input clk;
  input rst;
  output [7:0] fsm_output;
  reg [7:0] fsm_output;
  input Shift_Accum_Loop_C_5_tr0;


  // FSM State Type Declaration for fir_core_core_fsm_1
  parameter
    main_C_0 = 3'd0,
    Shift_Accum_Loop_C_0 = 3'd1,
    Shift_Accum_Loop_C_1 = 3'd2,
    Shift_Accum_Loop_C_2 = 3'd3,
    Shift_Accum_Loop_C_3 = 3'd4,
    Shift_Accum_Loop_C_4 = 3'd5,
    Shift_Accum_Loop_C_5 = 3'd6,
    main_C_1 = 3'd7;

  reg [2:0] state_var;
  reg [2:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : fir_core_core_fsm_1
    case (state_var)
      Shift_Accum_Loop_C_0 : begin
        fsm_output = 8'b00000010;
        state_var_NS = Shift_Accum_Loop_C_1;
      end
      Shift_Accum_Loop_C_1 : begin
        fsm_output = 8'b00000100;
        state_var_NS = Shift_Accum_Loop_C_2;
      end
      Shift_Accum_Loop_C_2 : begin
        fsm_output = 8'b00001000;
        state_var_NS = Shift_Accum_Loop_C_3;
      end
      Shift_Accum_Loop_C_3 : begin
        fsm_output = 8'b00010000;
        state_var_NS = Shift_Accum_Loop_C_4;
      end
      Shift_Accum_Loop_C_4 : begin
        fsm_output = 8'b00100000;
        state_var_NS = Shift_Accum_Loop_C_5;
      end
      Shift_Accum_Loop_C_5 : begin
        fsm_output = 8'b01000000;
        if ( Shift_Accum_Loop_C_5_tr0 ) begin
          state_var_NS = main_C_1;
        end
        else begin
          state_var_NS = Shift_Accum_Loop_C_0;
        end
      end
      main_C_1 : begin
        fsm_output = 8'b10000000;
        state_var_NS = main_C_0;
      end
      // main_C_0
      default : begin
        fsm_output = 8'b00000001;
        state_var_NS = Shift_Accum_Loop_C_0;
      end
    endcase
  end

  always @(posedge clk) begin
    if ( rst ) begin
      state_var <= main_C_0;
    end
    else begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    fir_core
// ------------------------------------------------------------------


module fir_core (
  clk, rst, y_rsc_dat, y_triosy_lz, x_rsc_dat, x_triosy_lz
);
  input clk;
  input rst;
  output [15:0] y_rsc_dat;
  output y_triosy_lz;
  input [7:0] x_rsc_dat;
  output x_triosy_lz;


  // Interconnect Declarations
  wire [7:0] x_rsci_idat;
  wire [7:0] fsm_output;
  wire or_tmp_13;
  wire or_tmp_16;
  reg i_3_sva;
  reg reg_x_triosy_obj_ld_cse;
  reg y_rsci_idat_rsp_0;
  reg [14:0] y_rsci_idat_rsp_1;
  wire reg_y_nor_ssc;
  reg [7:0] shift_reg_4_lpi_2;
  reg [7:0] shift_reg_3_lpi_2;
  reg [7:0] shift_reg_11_lpi_2;
  reg [7:0] shift_reg_2_lpi_2;
  reg [7:0] shift_reg_10_lpi_2;
  reg [7:0] shift_reg_9_lpi_2;
  reg [7:0] shift_reg_1_lpi_2;
  reg [7:0] shift_reg_0_lpi_2;
  reg [7:0] shift_reg_8_lpi_2;
  reg [7:0] shift_reg_7_lpi_2;
  reg [7:0] shift_reg_6_lpi_2;
  reg [7:0] shift_reg_5_lpi_2;
  reg [7:0] x_sva;
  reg acc_1_0_sva;
  wire [15:0] acc_6_sva_mx0w0;
  wire [17:0] nl_acc_6_sva_mx0w0;
  wire acc_6_sva_mx0c1;
  wire [7:0] Shift_Accum_Loop_3_else_Shift_Accum_Loop_else_slc_shift_reg_8_7_0_1_cse_sva_mx0;
  reg acc_6_sva_15;
  reg [14:0] acc_6_sva_14_0;
  wire or_cse;

  wire Shift_Accum_Loop_else_mux_1_nl;
  wire nor_nl;
  wire[12:0] Shift_Accum_Loop_acc_5_nl;
  wire[13:0] nl_Shift_Accum_Loop_acc_5_nl;
  wire[12:0] Shift_Accum_Loop_1_mul_nl;
  wire[7:0] shift_reg_static_init_else_mux_11_nl;
  wire[8:0] Shift_Accum_Loop_acc_8_nl;
  wire[9:0] nl_Shift_Accum_Loop_acc_8_nl;
  wire[12:0] Shift_Accum_Loop_5_mul_nl;
  wire[7:0] Shift_Accum_Loop_mux_2_nl;
  wire[14:0] and_67_nl;
  wire[14:0] Shift_Accum_Loop_acc_3_nl;
  wire[15:0] nl_Shift_Accum_Loop_acc_3_nl;
  wire[12:0] Shift_Accum_Loop_acc_7_nl;
  wire[13:0] nl_Shift_Accum_Loop_acc_7_nl;
  wire[7:0] Shift_Accum_Loop_acc_9_nl;
  wire[8:0] nl_Shift_Accum_Loop_acc_9_nl;
  wire acc_not_1_nl;
  wire mux_3_nl;
  wire mux_2_nl;
  wire or_32_nl;
  wire mux_1_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [15:0] nl_y_rsci_idat;
  assign nl_y_rsci_idat = {y_rsci_idat_rsp_0 , y_rsci_idat_rsp_1};
  wire  nl_fir_core_core_fsm_inst_Shift_Accum_Loop_C_5_tr0;
  assign nl_fir_core_core_fsm_inst_Shift_Accum_Loop_C_5_tr0 = ~ i_3_sva;
  ccs_out_v1 #(//.rscid(32'sd1),
  .width(32'sd16)) y_rsci (
      .idat(nl_y_rsci_idat[15:0]),
      .dat(y_rsc_dat)
    );
  ccs_in_v1 #(//.rscid(32'sd2),
  .width(32'sd8)) x_rsci (
      .dat(x_rsc_dat),
      .idat(x_rsci_idat)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) y_triosy_obj (
      .ld(reg_x_triosy_obj_ld_cse),
      .lz(y_triosy_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) x_triosy_obj (
      .ld(reg_x_triosy_obj_ld_cse),
      .lz(x_triosy_lz)
    );
  fir_core_core_fsm fir_core_core_fsm_inst (
      .clk(clk),
      .rst(rst),
      .fsm_output(fsm_output),
      .Shift_Accum_Loop_C_5_tr0(nl_fir_core_core_fsm_inst_Shift_Accum_Loop_C_5_tr0)
    );
  assign or_cse = (fsm_output[7]) | (fsm_output[0]);
  assign shift_reg_static_init_else_mux_11_nl = MUX_v_8_2_2(shift_reg_3_lpi_2, shift_reg_11_lpi_2,
      i_3_sva);
  assign Shift_Accum_Loop_1_mul_nl = shift_reg_static_init_else_mux_11_nl * ({(~
      i_3_sva) , 1'b0 , (~ i_3_sva) , 1'b0 , i_3_sva});
  assign nl_Shift_Accum_Loop_acc_8_nl = conv_u2u_8_9(Shift_Accum_Loop_3_else_Shift_Accum_Loop_else_slc_shift_reg_8_7_0_1_cse_sva_mx0)
      + conv_u2u_6_9(Shift_Accum_Loop_3_else_Shift_Accum_Loop_else_slc_shift_reg_8_7_0_1_cse_sva_mx0[7:2]);
  assign Shift_Accum_Loop_acc_8_nl = nl_Shift_Accum_Loop_acc_8_nl[8:0];
  assign nl_Shift_Accum_Loop_acc_5_nl = Shift_Accum_Loop_1_mul_nl + conv_u2u_12_13({Shift_Accum_Loop_acc_8_nl
      , (Shift_Accum_Loop_3_else_Shift_Accum_Loop_else_slc_shift_reg_8_7_0_1_cse_sva_mx0[1:0])
      , 1'b0});
  assign Shift_Accum_Loop_acc_5_nl = nl_Shift_Accum_Loop_acc_5_nl[12:0];
  assign Shift_Accum_Loop_mux_2_nl = MUX_v_8_2_2(x_sva, shift_reg_7_lpi_2, i_3_sva);
  assign Shift_Accum_Loop_5_mul_nl = Shift_Accum_Loop_mux_2_nl * ({i_3_sva , 1'b0
      , i_3_sva , 1'b0 , (~ i_3_sva)});
  assign nl_acc_6_sva_mx0w0 = ({acc_6_sva_14_0 , acc_1_0_sva}) + conv_u2u_13_16(Shift_Accum_Loop_acc_5_nl)
      + conv_u2u_13_16(Shift_Accum_Loop_5_mul_nl);
  assign acc_6_sva_mx0w0 = nl_acc_6_sva_mx0w0[15:0];
  assign Shift_Accum_Loop_3_else_Shift_Accum_Loop_else_slc_shift_reg_8_7_0_1_cse_sva_mx0
      = MUX_v_8_2_2(shift_reg_1_lpi_2, shift_reg_9_lpi_2, i_3_sva);
  assign or_tmp_13 = (~ (fsm_output[1])) | i_3_sva;
  assign or_tmp_16 = ~((fsm_output[1]) & i_3_sva);
  assign acc_6_sva_mx0c1 = (i_3_sva & (~ (fsm_output[7]))) | (fsm_output[6]) | (fsm_output[0]);
  assign reg_y_nor_ssc = ~((~ (fsm_output[6])) | i_3_sva);
  always @(posedge clk) begin
    if ( rst ) begin
      i_3_sva <= 1'b0;
    end
    else if ( (fsm_output[6]) | (fsm_output[0]) ) begin
      i_3_sva <= ~ (fsm_output[6]);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_sva <= 8'b00000000;
    end
    else if ( or_cse ) begin
      x_sva <= x_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      acc_1_0_sva <= 1'b0;
      reg_x_triosy_obj_ld_cse <= 1'b0;
    end
    else begin
      acc_1_0_sva <= Shift_Accum_Loop_else_mux_1_nl & (~ or_cse);
      reg_x_triosy_obj_ld_cse <= (~ i_3_sva) & (fsm_output[6]);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      shift_reg_1_lpi_2 <= 8'b00000000;
    end
    else if ( ~ or_tmp_13 ) begin
      shift_reg_1_lpi_2 <= shift_reg_0_lpi_2;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      shift_reg_3_lpi_2 <= 8'b00000000;
    end
    else if ( ~ or_tmp_13 ) begin
      shift_reg_3_lpi_2 <= shift_reg_2_lpi_2;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      shift_reg_5_lpi_2 <= 8'b00000000;
    end
    else if ( ~ or_tmp_16 ) begin
      shift_reg_5_lpi_2 <= shift_reg_4_lpi_2;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      shift_reg_7_lpi_2 <= 8'b00000000;
    end
    else if ( ~ or_tmp_16 ) begin
      shift_reg_7_lpi_2 <= shift_reg_6_lpi_2;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      shift_reg_9_lpi_2 <= 8'b00000000;
    end
    else if ( ~ or_tmp_16 ) begin
      shift_reg_9_lpi_2 <= shift_reg_8_lpi_2;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      shift_reg_11_lpi_2 <= 8'b00000000;
    end
    else if ( ~ or_tmp_16 ) begin
      shift_reg_11_lpi_2 <= shift_reg_10_lpi_2;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      shift_reg_0_lpi_2 <= 8'b00000000;
    end
    else if ( ~ or_tmp_13 ) begin
      shift_reg_0_lpi_2 <= x_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      shift_reg_2_lpi_2 <= 8'b00000000;
    end
    else if ( ~ or_tmp_13 ) begin
      shift_reg_2_lpi_2 <= shift_reg_1_lpi_2;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      shift_reg_6_lpi_2 <= 8'b00000000;
    end
    else if ( ~ or_tmp_16 ) begin
      shift_reg_6_lpi_2 <= shift_reg_5_lpi_2;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      shift_reg_8_lpi_2 <= 8'b00000000;
    end
    else if ( ~ or_tmp_16 ) begin
      shift_reg_8_lpi_2 <= shift_reg_7_lpi_2;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      shift_reg_10_lpi_2 <= 8'b00000000;
    end
    else if ( ~ or_tmp_16 ) begin
      shift_reg_10_lpi_2 <= shift_reg_9_lpi_2;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      shift_reg_4_lpi_2 <= 8'b00000000;
    end
    else if ( fsm_output[1] ) begin
      shift_reg_4_lpi_2 <= shift_reg_3_lpi_2;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      y_rsci_idat_rsp_0 <= 1'b0;
      y_rsci_idat_rsp_1 <= 15'b000000000000000;
    end
    else if ( reg_y_nor_ssc ) begin
      y_rsci_idat_rsp_0 <= acc_6_sva_15;
      y_rsci_idat_rsp_1 <= acc_6_sva_14_0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      acc_6_sva_15 <= 1'b0;
    end
    else if ( ((~ i_3_sva) & (fsm_output[1])) | acc_6_sva_mx0c1 ) begin
      acc_6_sva_15 <= acc_6_sva_mx0w0[15];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      acc_6_sva_14_0 <= 15'b000000000000000;
    end
    else if ( mux_3_nl | (fsm_output[0]) ) begin
      acc_6_sva_14_0 <= MUX_v_15_2_2((acc_6_sva_mx0w0[14:0]), and_67_nl, acc_6_sva_mx0c1);
    end
  end
  assign nor_nl = ~((fsm_output[1]) | (fsm_output[7]) | (fsm_output[0]));
  assign Shift_Accum_Loop_else_mux_1_nl = MUX_s_1_2_2((acc_6_sva_mx0w0[0]), acc_1_0_sva,
      nor_nl);
  assign nl_Shift_Accum_Loop_acc_9_nl = conv_u2s_5_8(shift_reg_5_lpi_2[7:3]) + (~
      shift_reg_5_lpi_2);
  assign Shift_Accum_Loop_acc_9_nl = nl_Shift_Accum_Loop_acc_9_nl[7:0];
  assign nl_Shift_Accum_Loop_acc_7_nl = ({shift_reg_5_lpi_2 , 5'b01000}) + conv_s2u_12_13({1'b1
      , Shift_Accum_Loop_acc_9_nl , (shift_reg_5_lpi_2[2:0])});
  assign Shift_Accum_Loop_acc_7_nl = nl_Shift_Accum_Loop_acc_7_nl[12:0];
  assign nl_Shift_Accum_Loop_acc_3_nl = conv_u2u_13_15(Shift_Accum_Loop_acc_7_nl)
      + (acc_6_sva_mx0w0[15:1]);
  assign Shift_Accum_Loop_acc_3_nl = nl_Shift_Accum_Loop_acc_3_nl[14:0];
  assign acc_not_1_nl = ~ or_cse;
  assign and_67_nl = MUX_v_15_2_2(15'b000000000000000, Shift_Accum_Loop_acc_3_nl,
      acc_not_1_nl);
  assign or_32_nl = (fsm_output[1]) | (fsm_output[6]);
  assign mux_2_nl = MUX_s_1_2_2((fsm_output[1]), or_32_nl, fsm_output[7]);
  assign mux_1_nl = MUX_s_1_2_2((fsm_output[1]), (fsm_output[6]), fsm_output[7]);
  assign mux_3_nl = MUX_s_1_2_2(mux_2_nl, mux_1_nl, i_3_sva);

  function automatic  MUX_s_1_2_2;
    input  input_0;
    input  input_1;
    input  sel;
    reg  result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [14:0] MUX_v_15_2_2;
    input [14:0] input_0;
    input [14:0] input_1;
    input  sel;
    reg [14:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_15_2_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input  sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction


  function automatic [12:0] conv_s2u_12_13 ;
    input [11:0]  vector ;
  begin
    conv_s2u_12_13 = {vector[11], vector};
  end
  endfunction


  function automatic [7:0] conv_u2s_5_8 ;
    input [4:0]  vector ;
  begin
    conv_u2s_5_8 = {{3{1'b0}}, vector};
  end
  endfunction


  function automatic [8:0] conv_u2u_6_9 ;
    input [5:0]  vector ;
  begin
    conv_u2u_6_9 = {{3{1'b0}}, vector};
  end
  endfunction


  function automatic [8:0] conv_u2u_8_9 ;
    input [7:0]  vector ;
  begin
    conv_u2u_8_9 = {1'b0, vector};
  end
  endfunction


  function automatic [12:0] conv_u2u_12_13 ;
    input [11:0]  vector ;
  begin
    conv_u2u_12_13 = {1'b0, vector};
  end
  endfunction


  function automatic [14:0] conv_u2u_13_15 ;
    input [12:0]  vector ;
  begin
    conv_u2u_13_15 = {{2{1'b0}}, vector};
  end
  endfunction


  function automatic [15:0] conv_u2u_13_16 ;
    input [12:0]  vector ;
  begin
    conv_u2u_13_16 = {{3{1'b0}}, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    fir
// ------------------------------------------------------------------


module fir (
  clk, rst, y_rsc_dat, y_triosy_lz, x_rsc_dat, x_triosy_lz
);
  input clk;
  input rst;
  output [15:0] y_rsc_dat;
  output y_triosy_lz;
  input [7:0] x_rsc_dat;
  output x_triosy_lz;



  // Interconnect Declarations for Component Instantiations 
  fir_core fir_core_inst (
      .clk(clk),
      .rst(rst),
      .y_rsc_dat(y_rsc_dat),
      .y_triosy_lz(y_triosy_lz),
      .x_rsc_dat(x_rsc_dat),
      .x_triosy_lz(x_triosy_lz)
    );
endmodule


